`timescale 1ps / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:21:52 02/02/2021 
// Design Name: 
// Module Name:    top_riscv 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module top_riscv_pl(top_dmemrw,top_dmem_data,top_dmem_addr,top_dmem_out,top_imem_addr,top_imem_inst,clk,rst
    );
	 
///////////////////////////////////////////////////////////////////////////////////Ports Declaration section///////////////////////////////////////////////////////////
/////////////////////////////////////////Data memory ports///////////////////////////////////
	 input  [31:0] top_dmem_out                ;
	 output [31:0] top_dmem_data,top_dmem_addr ;
	 output        top_dmemrw                  ;
//////////////////////////////////////////////////////////////////////////////////////////////
	 
/////////////////////////////////////Instruction memory ports/////////////////////////////////
	 input   [31:0] top_imem_inst              ;
	 output  [31:0] top_imem_addr              ;
//////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////Global ports///////////////////////////////// //////////
	input           clk,rst                    ;
//////////////////////////////////////////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////End of section/////////////////////////////////////////////////////////////////////


///////////////////////////////////////////////////////////////////////////////////Internal regs and wires section////////////////////////////////////////////////////
	wire [2:0]  dp_cl_immsel	                    ;
	wire [1:0]  dp_cl_wbsel                        ;
	wire        dp_cl_pcsel,dp_cl_regwen           ;
	wire			dp_cl_brun,dp_cl_breq,dp_cl_brlt   ;
	wire        dp_cl_asel,dp_cl_bsel              ;
	wire [3:0]  dp_cl_alusel                       ;
	wire [31:0] dp_cl_instr_pl							  ;
	wire        dp_cl_dmemrw							  ;
	wire [31:0] wb_reg_out,regw_reg_out				  ;
///////////////////////////////////////////////////////////////////////////////////End of section/////////////////////////////////////////////////////////////////////


///////////////////////////////////////////////////////////////////////////////////combinational section////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////////End of section/////////////////////////////////////////////////////////////////////
assign top_dmemrw=wb_reg_out[2];

///////////////////////////////////////////////////////////////////////////////////Components section////////////////////////////////////////////////////
top_dp_pl       dp (.dp_rst(rst) , .dp_clk (clk) , .dp_pcsel(dp_cl_pcsel)  , .dp_immsel(dp_cl_immsel) , .dp_regwen(regw_reg_out[0]) , .dp_datab(top_dmem_data)       ,  //DP instance
					  .dp_brun(dp_cl_brun) , .dp_brlt(dp_cl_brlt) , .dp_breq(dp_cl_breq) , .dp_bsel(dp_cl_bsel) , .dp_asel(dp_cl_asel) , .dp_alusel(dp_cl_alusel)   ,
					  .dp_wbsel(wb_reg_out[1:0]) , .dp_dmem_out(top_dmem_out) , .dp_imem_inst(top_imem_inst) , .dp_pc_next(top_imem_addr) , .dp_alu_out(top_dmem_addr),.pl_inst(dp_cl_instr_pl)) ;
					  
reg_mod			 wb_reg(.data_in({28'b0,dp_cl_regwen,dp_cl_dmemrw,dp_cl_wbsel}) ,.data_out(wb_reg_out) ,.clk(clk),.rst(rst));

reg_mod         regw_reg(.data_in({31'b0,wb_reg_out[3]}),.data_out(regw_reg_out) ,.clk(clk),.rst(rst));
					  
Control_Unit cl (.instr(dp_cl_instr_pl) , .breq(dp_cl_breq) , .brlt(dp_cl_brlt) , .pc_sel(dp_cl_pcsel) , .a_sel(dp_cl_asel) , .b_sel(dp_cl_bsel)                 ,  //Control logic instance
					  .mem_write_en(dp_cl_dmemrw) , .reg_file_wr_en(dp_cl_regwen) , .alu_sel(dp_cl_alusel) , .wb_sel(dp_cl_wbsel) , .imm_sel(dp_cl_immsel)            ,
					  .pr_un(dp_cl_brun))                                                                                                                           ;

///////////////////////////////////////////////////////////////////////////////////End of section/////////////////////////////////////////////////////////////////////
endmodule
